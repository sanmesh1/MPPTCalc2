* C:\Users\sanme_000\Documents\Visual Studio 2015\Projects\VideoRental2\VideoRental2\Content\OtherFile\RC2.asc
V1 N001 0 5
C1 N002 0 1m
R1 N001 N002 5
.ic v(n002) = 0
.tran 25m
.backanno
.end
